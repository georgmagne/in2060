library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.numeric_std.all;

  -- Denne kildekoden har lagt inn 2 skrivefeil.
  -- Skriv koden selv, og kommenter feilene der du finner dem.

entity MAC is
    generic (width: integer := 8);
    port(
        clk, reset  : in STD_LOGIC; -- Første feil, mangler semikolon
        MLS_select  : in STD_LOGIC;
        Rn, Rm, Ra  : in STD_LOGIC_VECTOR(width-1 downto 0);
        Rd          : out STD_LOGIC_VECTOR(width-1 downto 0)
    );
    end;

architecture behavioral of MAC is
    signal mul1, mul2, add1, buffRa 	: UNSIGNED(width-1 downto 0);     -- Lagt til buffRa, som buffer til Ra.
    signal add2, sum, buffProd        : UNSIGNED(width*2-1 downto 0);   -- Lagt til buffProd, som buffer til produktet Rm*Rn.

    begin
      process(clk, reset)

      begin
        if reset = '1' then
          Rd <= (others => '0');                  -- asynkron reset.
          buffProd <= (others => '0');            -- Resetter bufferene
          buffRa <= (others => '0');

      elsif rising_edge(clk) then                 -- Skjer på positiv klokkeflanke.
        buffProd <= add2;                         -- buffProd settes til produktet til Rn*Rm
        buffRa <= add1;                           -- buddRa settes til verdien Ra har
        
        Rd <= STD_LOGIC_VECTOR(sum(width-1 downto 0)); -- Ta vare på LSB. -- Andre feil, sum var sm.
      end if;

    end process;

    -- Concurrent statements
    -- Skjer utenfor prosess, uavhening av klokkeflanker.

    mul1 <= UNSIGNED(Rn);
    mul2 <= UNSIGNED(Rm);
    add1 <= UNSIGNED(Ra);
    add2 <= mul1*mul2;
    sum <= buffRa + buffProd;    -- Ender sum til å være summen av bufferene til Ra og Rn*Rm.

  end architecture;
